Parallel2Serial_32bits_inst : Parallel2Serial_32bits PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		load	 => load_sig,
		shiftout	 => shiftout_sig
	);
