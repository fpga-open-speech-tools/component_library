Serial2Parallel_32bits_inst : Serial2Parallel_32bits PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		q	 => q_sig
	);
