library IEEE;
use IEEE.std_logic_1164.all;

package ad1939 is

  constant word_length : integer := 24; 
  constant fraction_length : integer := 23;

end package;